// HPSWrapper.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module HPSWrapper (
		input  wire [29:0] ddr_read_address,                 //        ddr_read.address
		input  wire [7:0]  ddr_read_burstcount,              //                .burstcount
		output wire        ddr_read_waitrequest,             //                .waitrequest
		output wire [31:0] ddr_read_readdata,                //                .readdata
		output wire        ddr_read_readdatavalid,           //                .readdatavalid
		input  wire        ddr_read_read,                    //                .read
		input  wire        ddr_read_clock_clk,               //  ddr_read_clock.clk
		output wire        ddr_read_reset_reset,             //  ddr_read_reset.reset
		input  wire [29:0] ddr_write_address,                //       ddr_write.address
		input  wire [7:0]  ddr_write_burstcount,             //                .burstcount
		output wire        ddr_write_waitrequest,            //                .waitrequest
		input  wire [31:0] ddr_write_writedata,              //                .writedata
		input  wire [3:0]  ddr_write_byteenable,             //                .byteenable
		input  wire        ddr_write_write,                  //                .write
		input  wire        ddr_write_clock_clk,              // ddr_write_clock.clk
		output wire        ddr_write_reset_reset,            // ddr_write_reset.reset
		input  wire [16:0] handshake_in_port,                //       handshake.in_port
		output wire [16:0] handshake_out_port,               //                .out_port
		output wire        hps_avmm_master_chipselect,       // hps_avmm_master.chipselect
		output wire        hps_avmm_master_read,             //                .read
		input  wire [31:0] hps_avmm_master_readdata,         //                .readdata
		output wire [31:0] hps_avmm_master_writedata,        //                .writedata
		output wire        hps_avmm_master_write,            //                .write
		output wire [3:0]  hps_avmm_master_byteenable,       //                .byteenable
		output wire [13:0] hps_avmm_master_address,          //                .address
		inout  wire        hps_io_hps_io_sdio_inst_CMD,      //          hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,       //                .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,       //                .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,      //                .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,       //                .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,       //                .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,      //                .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,      //                .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,   //                .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,   //                .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,   //                .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO49, //                .hps_io_gpio_inst_LOANIO49
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO50, //                .hps_io_gpio_inst_LOANIO50
		output wire        lt24_cmd_ready,                   //        lt24_cmd.ready
		input  wire [7:0]  lt24_cmd_data,                    //                .data
		input  wire        lt24_cmd_write,                   //                .write
		input  wire        lt24_cmd_done,                    //                .done
		output wire        lt24_data_ready,                  //       lt24_data.ready
		input  wire [15:0] lt24_data_data,                   //                .data
		input  wire        lt24_data_write,                  //                .write
		input  wire [7:0]  lt24_data_xAddr,                  //                .xAddr
		input  wire [8:0]  lt24_data_yAddr,                  //                .yAddr
		output wire        lt24_display_cs_n,                //    lt24_display.cs_n
		output wire        lt24_display_rs,                  //                .rs
		output wire        lt24_display_rd_n,                //                .rd_n
		output wire        lt24_display_wr_n,                //                .wr_n
		output wire [15:0] lt24_display_data,                //                .data
		output wire        lt24_display_on,                  //                .on
		output wire        lt24_display_rst_n,               //                .rst_n
		input  wire        lt24_mode_raw,                    //       lt24_mode.raw
		output wire [14:0] memory_mem_a,                     //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //                .mem_ba
		output wire        memory_mem_ck,                    //                .mem_ck
		output wire        memory_mem_ck_n,                  //                .mem_ck_n
		output wire        memory_mem_cke,                   //                .mem_cke
		output wire        memory_mem_cs_n,                  //                .mem_cs_n
		output wire        memory_mem_ras_n,                 //                .mem_ras_n
		output wire        memory_mem_cas_n,                 //                .mem_cas_n
		output wire        memory_mem_we_n,                  //                .mem_we_n
		output wire        memory_mem_reset_n,               //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                    //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                   //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                 //                .mem_dqs_n
		output wire        memory_mem_odt,                   //                .mem_odt
		output wire [3:0]  memory_mem_dm,                    //                .mem_dm
		input  wire        memory_oct_rzqin,                 //                .oct_rzqin
		output wire        usb_uart_rx,                      //        usb_uart.rx
		input  wire        usb_uart_tx,                      //                .tx
		input  wire        user_clock_clk,                   //      user_clock.clk
		output wire        user_reset_reset                  //      user_reset.reset
	);

	wire         reset_width_overflow_overflow;                      // reset_width:overflow -> hps_reset:sigIn
	wire  [66:0] arm_hps_h2f_loan_io_in;                             // arm_hps:h2f_loan_in -> usb_uart:loan_io_in
	wire  [66:0] usb_uart_loan_io_oe;                                // usb_uart:loan_io_oe -> arm_hps:h2f_loan_oe
	wire  [66:0] usb_uart_loan_io_out;                               // usb_uart:loan_io_out -> arm_hps:h2f_loan_out
	wire         arm_hps_h2f_reset_reset;                            // arm_hps:h2f_rst_n -> [reset50mhz:reset_in0, rst_controller_001:reset_in0]
	wire         power_on_reset_reset_reset;                         // power_on_reset:reset -> [hps_reset:reset, reset50mhz:reset_in2, reset_width:reset]
	wire         hps_reset_reset_reset;                              // hps_reset:sigOut -> [arm_hps:f2h_cold_rst_req_n, reset50mhz:reset_in1]
	wire         hpsinitreset_user_reset_reset;                      // hpsInitReset:user_reset -> [ddr_read_rst:reset_in0, ddr_write_rst:reset_in0, lt24_fpga:globalReset]
	wire   [1:0] arm_hps_h2f_axi_master_awburst;                     // arm_hps:h2f_AWBURST -> mm_interconnect_0:arm_hps_h2f_axi_master_awburst
	wire   [3:0] arm_hps_h2f_axi_master_arlen;                       // arm_hps:h2f_ARLEN -> mm_interconnect_0:arm_hps_h2f_axi_master_arlen
	wire   [3:0] arm_hps_h2f_axi_master_wstrb;                       // arm_hps:h2f_WSTRB -> mm_interconnect_0:arm_hps_h2f_axi_master_wstrb
	wire         arm_hps_h2f_axi_master_wready;                      // mm_interconnect_0:arm_hps_h2f_axi_master_wready -> arm_hps:h2f_WREADY
	wire  [11:0] arm_hps_h2f_axi_master_rid;                         // mm_interconnect_0:arm_hps_h2f_axi_master_rid -> arm_hps:h2f_RID
	wire         arm_hps_h2f_axi_master_rready;                      // arm_hps:h2f_RREADY -> mm_interconnect_0:arm_hps_h2f_axi_master_rready
	wire   [3:0] arm_hps_h2f_axi_master_awlen;                       // arm_hps:h2f_AWLEN -> mm_interconnect_0:arm_hps_h2f_axi_master_awlen
	wire  [11:0] arm_hps_h2f_axi_master_wid;                         // arm_hps:h2f_WID -> mm_interconnect_0:arm_hps_h2f_axi_master_wid
	wire   [3:0] arm_hps_h2f_axi_master_arcache;                     // arm_hps:h2f_ARCACHE -> mm_interconnect_0:arm_hps_h2f_axi_master_arcache
	wire         arm_hps_h2f_axi_master_wvalid;                      // arm_hps:h2f_WVALID -> mm_interconnect_0:arm_hps_h2f_axi_master_wvalid
	wire  [29:0] arm_hps_h2f_axi_master_araddr;                      // arm_hps:h2f_ARADDR -> mm_interconnect_0:arm_hps_h2f_axi_master_araddr
	wire   [2:0] arm_hps_h2f_axi_master_arprot;                      // arm_hps:h2f_ARPROT -> mm_interconnect_0:arm_hps_h2f_axi_master_arprot
	wire   [2:0] arm_hps_h2f_axi_master_awprot;                      // arm_hps:h2f_AWPROT -> mm_interconnect_0:arm_hps_h2f_axi_master_awprot
	wire  [31:0] arm_hps_h2f_axi_master_wdata;                       // arm_hps:h2f_WDATA -> mm_interconnect_0:arm_hps_h2f_axi_master_wdata
	wire         arm_hps_h2f_axi_master_arvalid;                     // arm_hps:h2f_ARVALID -> mm_interconnect_0:arm_hps_h2f_axi_master_arvalid
	wire   [3:0] arm_hps_h2f_axi_master_awcache;                     // arm_hps:h2f_AWCACHE -> mm_interconnect_0:arm_hps_h2f_axi_master_awcache
	wire  [11:0] arm_hps_h2f_axi_master_arid;                        // arm_hps:h2f_ARID -> mm_interconnect_0:arm_hps_h2f_axi_master_arid
	wire   [1:0] arm_hps_h2f_axi_master_arlock;                      // arm_hps:h2f_ARLOCK -> mm_interconnect_0:arm_hps_h2f_axi_master_arlock
	wire   [1:0] arm_hps_h2f_axi_master_awlock;                      // arm_hps:h2f_AWLOCK -> mm_interconnect_0:arm_hps_h2f_axi_master_awlock
	wire  [29:0] arm_hps_h2f_axi_master_awaddr;                      // arm_hps:h2f_AWADDR -> mm_interconnect_0:arm_hps_h2f_axi_master_awaddr
	wire   [1:0] arm_hps_h2f_axi_master_bresp;                       // mm_interconnect_0:arm_hps_h2f_axi_master_bresp -> arm_hps:h2f_BRESP
	wire         arm_hps_h2f_axi_master_arready;                     // mm_interconnect_0:arm_hps_h2f_axi_master_arready -> arm_hps:h2f_ARREADY
	wire  [31:0] arm_hps_h2f_axi_master_rdata;                       // mm_interconnect_0:arm_hps_h2f_axi_master_rdata -> arm_hps:h2f_RDATA
	wire         arm_hps_h2f_axi_master_awready;                     // mm_interconnect_0:arm_hps_h2f_axi_master_awready -> arm_hps:h2f_AWREADY
	wire   [1:0] arm_hps_h2f_axi_master_arburst;                     // arm_hps:h2f_ARBURST -> mm_interconnect_0:arm_hps_h2f_axi_master_arburst
	wire   [2:0] arm_hps_h2f_axi_master_arsize;                      // arm_hps:h2f_ARSIZE -> mm_interconnect_0:arm_hps_h2f_axi_master_arsize
	wire         arm_hps_h2f_axi_master_bready;                      // arm_hps:h2f_BREADY -> mm_interconnect_0:arm_hps_h2f_axi_master_bready
	wire         arm_hps_h2f_axi_master_rlast;                       // mm_interconnect_0:arm_hps_h2f_axi_master_rlast -> arm_hps:h2f_RLAST
	wire         arm_hps_h2f_axi_master_wlast;                       // arm_hps:h2f_WLAST -> mm_interconnect_0:arm_hps_h2f_axi_master_wlast
	wire   [1:0] arm_hps_h2f_axi_master_rresp;                       // mm_interconnect_0:arm_hps_h2f_axi_master_rresp -> arm_hps:h2f_RRESP
	wire  [11:0] arm_hps_h2f_axi_master_awid;                        // arm_hps:h2f_AWID -> mm_interconnect_0:arm_hps_h2f_axi_master_awid
	wire  [11:0] arm_hps_h2f_axi_master_bid;                         // mm_interconnect_0:arm_hps_h2f_axi_master_bid -> arm_hps:h2f_BID
	wire         arm_hps_h2f_axi_master_bvalid;                      // mm_interconnect_0:arm_hps_h2f_axi_master_bvalid -> arm_hps:h2f_BVALID
	wire   [2:0] arm_hps_h2f_axi_master_awsize;                      // arm_hps:h2f_AWSIZE -> mm_interconnect_0:arm_hps_h2f_axi_master_awsize
	wire         arm_hps_h2f_axi_master_awvalid;                     // arm_hps:h2f_AWVALID -> mm_interconnect_0:arm_hps_h2f_axi_master_awvalid
	wire         arm_hps_h2f_axi_master_rvalid;                      // mm_interconnect_0:arm_hps_h2f_axi_master_rvalid -> arm_hps:h2f_RVALID
	wire         mm_interconnect_0_baremetal_s1_chipselect;          // mm_interconnect_0:baremetal_s1_chipselect -> baremetal:chipselect
	wire  [31:0] mm_interconnect_0_baremetal_s1_readdata;            // baremetal:readdata -> mm_interconnect_0:baremetal_s1_readdata
	wire         mm_interconnect_0_baremetal_s1_debugaccess;         // mm_interconnect_0:baremetal_s1_debugaccess -> baremetal:debugaccess
	wire  [13:0] mm_interconnect_0_baremetal_s1_address;             // mm_interconnect_0:baremetal_s1_address -> baremetal:address
	wire   [3:0] mm_interconnect_0_baremetal_s1_byteenable;          // mm_interconnect_0:baremetal_s1_byteenable -> baremetal:byteenable
	wire         mm_interconnect_0_baremetal_s1_write;               // mm_interconnect_0:baremetal_s1_write -> baremetal:write
	wire  [31:0] mm_interconnect_0_baremetal_s1_writedata;           // mm_interconnect_0:baremetal_s1_writedata -> baremetal:writedata
	wire         mm_interconnect_0_baremetal_s1_clken;               // mm_interconnect_0:baremetal_s1_clken -> baremetal:clken
	wire   [1:0] arm_hps_h2f_lw_axi_master_awburst;                  // arm_hps:h2f_lw_AWBURST -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awburst
	wire   [3:0] arm_hps_h2f_lw_axi_master_arlen;                    // arm_hps:h2f_lw_ARLEN -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arlen
	wire   [3:0] arm_hps_h2f_lw_axi_master_wstrb;                    // arm_hps:h2f_lw_WSTRB -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_wstrb
	wire         arm_hps_h2f_lw_axi_master_wready;                   // mm_interconnect_1:arm_hps_h2f_lw_axi_master_wready -> arm_hps:h2f_lw_WREADY
	wire  [11:0] arm_hps_h2f_lw_axi_master_rid;                      // mm_interconnect_1:arm_hps_h2f_lw_axi_master_rid -> arm_hps:h2f_lw_RID
	wire         arm_hps_h2f_lw_axi_master_rready;                   // arm_hps:h2f_lw_RREADY -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_rready
	wire   [3:0] arm_hps_h2f_lw_axi_master_awlen;                    // arm_hps:h2f_lw_AWLEN -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awlen
	wire  [11:0] arm_hps_h2f_lw_axi_master_wid;                      // arm_hps:h2f_lw_WID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_wid
	wire   [3:0] arm_hps_h2f_lw_axi_master_arcache;                  // arm_hps:h2f_lw_ARCACHE -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arcache
	wire         arm_hps_h2f_lw_axi_master_wvalid;                   // arm_hps:h2f_lw_WVALID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_hps_h2f_lw_axi_master_araddr;                   // arm_hps:h2f_lw_ARADDR -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_araddr
	wire   [2:0] arm_hps_h2f_lw_axi_master_arprot;                   // arm_hps:h2f_lw_ARPROT -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arprot
	wire   [2:0] arm_hps_h2f_lw_axi_master_awprot;                   // arm_hps:h2f_lw_AWPROT -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awprot
	wire  [31:0] arm_hps_h2f_lw_axi_master_wdata;                    // arm_hps:h2f_lw_WDATA -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_wdata
	wire         arm_hps_h2f_lw_axi_master_arvalid;                  // arm_hps:h2f_lw_ARVALID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_hps_h2f_lw_axi_master_awcache;                  // arm_hps:h2f_lw_AWCACHE -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awcache
	wire  [11:0] arm_hps_h2f_lw_axi_master_arid;                     // arm_hps:h2f_lw_ARID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arid
	wire   [1:0] arm_hps_h2f_lw_axi_master_arlock;                   // arm_hps:h2f_lw_ARLOCK -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arlock
	wire   [1:0] arm_hps_h2f_lw_axi_master_awlock;                   // arm_hps:h2f_lw_AWLOCK -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awlock
	wire  [20:0] arm_hps_h2f_lw_axi_master_awaddr;                   // arm_hps:h2f_lw_AWADDR -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_hps_h2f_lw_axi_master_bresp;                    // mm_interconnect_1:arm_hps_h2f_lw_axi_master_bresp -> arm_hps:h2f_lw_BRESP
	wire         arm_hps_h2f_lw_axi_master_arready;                  // mm_interconnect_1:arm_hps_h2f_lw_axi_master_arready -> arm_hps:h2f_lw_ARREADY
	wire  [31:0] arm_hps_h2f_lw_axi_master_rdata;                    // mm_interconnect_1:arm_hps_h2f_lw_axi_master_rdata -> arm_hps:h2f_lw_RDATA
	wire         arm_hps_h2f_lw_axi_master_awready;                  // mm_interconnect_1:arm_hps_h2f_lw_axi_master_awready -> arm_hps:h2f_lw_AWREADY
	wire   [1:0] arm_hps_h2f_lw_axi_master_arburst;                  // arm_hps:h2f_lw_ARBURST -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arburst
	wire   [2:0] arm_hps_h2f_lw_axi_master_arsize;                   // arm_hps:h2f_lw_ARSIZE -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_arsize
	wire         arm_hps_h2f_lw_axi_master_bready;                   // arm_hps:h2f_lw_BREADY -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_bready
	wire         arm_hps_h2f_lw_axi_master_rlast;                    // mm_interconnect_1:arm_hps_h2f_lw_axi_master_rlast -> arm_hps:h2f_lw_RLAST
	wire         arm_hps_h2f_lw_axi_master_wlast;                    // arm_hps:h2f_lw_WLAST -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_wlast
	wire   [1:0] arm_hps_h2f_lw_axi_master_rresp;                    // mm_interconnect_1:arm_hps_h2f_lw_axi_master_rresp -> arm_hps:h2f_lw_RRESP
	wire  [11:0] arm_hps_h2f_lw_axi_master_awid;                     // arm_hps:h2f_lw_AWID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awid
	wire  [11:0] arm_hps_h2f_lw_axi_master_bid;                      // mm_interconnect_1:arm_hps_h2f_lw_axi_master_bid -> arm_hps:h2f_lw_BID
	wire         arm_hps_h2f_lw_axi_master_bvalid;                   // mm_interconnect_1:arm_hps_h2f_lw_axi_master_bvalid -> arm_hps:h2f_lw_BVALID
	wire   [2:0] arm_hps_h2f_lw_axi_master_awsize;                   // arm_hps:h2f_lw_AWSIZE -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awsize
	wire         arm_hps_h2f_lw_axi_master_awvalid;                  // arm_hps:h2f_lw_AWVALID -> mm_interconnect_1:arm_hps_h2f_lw_axi_master_awvalid
	wire         arm_hps_h2f_lw_axi_master_rvalid;                   // mm_interconnect_1:arm_hps_h2f_lw_axi_master_rvalid -> arm_hps:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;     // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;      // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_handshake_s1_chipselect;          // mm_interconnect_1:handshake_s1_chipselect -> handshake:chipselect
	wire  [31:0] mm_interconnect_1_handshake_s1_readdata;            // handshake:readdata -> mm_interconnect_1:handshake_s1_readdata
	wire   [1:0] mm_interconnect_1_handshake_s1_address;             // mm_interconnect_1:handshake_s1_address -> handshake:address
	wire         mm_interconnect_1_handshake_s1_write;               // mm_interconnect_1:handshake_s1_write -> handshake:write_n
	wire  [31:0] mm_interconnect_1_handshake_s1_writedata;           // mm_interconnect_1:handshake_s1_writedata -> handshake:writedata
	wire         mm_interconnect_1_hps_avmm_master_slave_chipselect; // mm_interconnect_1:hps_avmm_master_slave_chipselect -> hps_avmm_master:slave_chip_sel
	wire  [31:0] mm_interconnect_1_hps_avmm_master_slave_readdata;   // hps_avmm_master:slave_readdata -> mm_interconnect_1:hps_avmm_master_slave_readdata
	wire  [13:0] mm_interconnect_1_hps_avmm_master_slave_address;    // mm_interconnect_1:hps_avmm_master_slave_address -> hps_avmm_master:slave_address
	wire         mm_interconnect_1_hps_avmm_master_slave_read;       // mm_interconnect_1:hps_avmm_master_slave_read -> hps_avmm_master:slave_read
	wire   [3:0] mm_interconnect_1_hps_avmm_master_slave_byteenable; // mm_interconnect_1:hps_avmm_master_slave_byteenable -> hps_avmm_master:slave_byte_en
	wire         mm_interconnect_1_hps_avmm_master_slave_write;      // mm_interconnect_1:hps_avmm_master_slave_write -> hps_avmm_master:slave_write
	wire  [31:0] mm_interconnect_1_hps_avmm_master_slave_writedata;  // mm_interconnect_1:hps_avmm_master_slave_writedata -> hps_avmm_master:slave_writedata
	wire         mm_interconnect_1_hpsinitreset_slave_chipselect;    // mm_interconnect_1:hpsInitReset_slave_chipselect -> hpsInitReset:chipsel
	wire         mm_interconnect_1_hpsinitreset_slave_write;         // mm_interconnect_1:hpsInitReset_slave_write -> hpsInitReset:write
	wire  [31:0] mm_interconnect_1_hpsinitreset_slave_writedata;     // mm_interconnect_1:hpsInitReset_slave_writedata -> hpsInitReset:writedata
	wire         irq_mapper_receiver0_irq;                           // handshake:irq -> irq_mapper:receiver0_irq
	wire  [31:0] arm_hps_f2h_irq0_irq;                               // irq_mapper:sender_irq -> arm_hps:f2h_irq_p0
	wire  [31:0] arm_hps_f2h_irq1_irq;                               // irq_mapper_001:sender_irq -> arm_hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [baremetal:reset, hpsInitReset:reset, mm_interconnect_0:baremetal_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:sysid_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [baremetal:reset_req, rst_translator:reset_req_in]
	wire         reset50mhz_reset_out_reset;                         // reset50mhz:reset_out -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> [mm_interconnect_0:arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:arm_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	HPSWrapper_arm_hps #(
		.F2S_Width (0),
		.S2F_Width (1)
	) arm_hps (
		.h2f_loan_in               (arm_hps_h2f_loan_io_in),            //        h2f_loan_io.in
		.h2f_loan_out              (usb_uart_loan_io_out),              //                   .out
		.h2f_loan_oe               (usb_uart_loan_io_oe),               //                   .oe
		.f2h_cold_rst_req_n        (hps_reset_reset_reset),             // f2h_cold_reset_req.reset_n
		.mem_a                     (memory_mem_a),                      //             memory.mem_a
		.mem_ba                    (memory_mem_ba),                     //                   .mem_ba
		.mem_ck                    (memory_mem_ck),                     //                   .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                   //                   .mem_ck_n
		.mem_cke                   (memory_mem_cke),                    //                   .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                   //                   .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                  //                   .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                  //                   .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                   //                   .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                //                   .mem_reset_n
		.mem_dq                    (memory_mem_dq),                     //                   .mem_dq
		.mem_dqs                   (memory_mem_dqs),                    //                   .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                  //                   .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                    //                   .mem_odt
		.mem_dm                    (memory_mem_dm),                     //                   .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                  //                   .oct_rzqin
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),       //             hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),        //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),        //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),       //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),        //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),        //                   .hps_io_sdio_inst_D3
		.hps_io_i2c0_inst_SDA      (hps_io_hps_io_i2c0_inst_SDA),       //                   .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_io_hps_io_i2c0_inst_SCL),       //                   .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO48   (hps_io_hps_io_gpio_inst_GPIO48),    //                   .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53   (hps_io_hps_io_gpio_inst_GPIO53),    //                   .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54   (hps_io_hps_io_gpio_inst_GPIO54),    //                   .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_LOANIO49 (hps_io_hps_io_gpio_inst_LOANIO49),  //                   .hps_io_gpio_inst_LOANIO49
		.hps_io_gpio_inst_LOANIO50 (hps_io_hps_io_gpio_inst_LOANIO50),  //                   .hps_io_gpio_inst_LOANIO50
		.h2f_rst_n                 (arm_hps_h2f_reset_reset),           //          h2f_reset.reset_n
		.f2h_sdram0_clk            (ddr_read_clock_clk),                //   f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS        (ddr_read_address),                  //    f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT     (ddr_read_burstcount),               //                   .burstcount
		.f2h_sdram0_WAITREQUEST    (ddr_read_waitrequest),              //                   .waitrequest
		.f2h_sdram0_READDATA       (ddr_read_readdata),                 //                   .readdata
		.f2h_sdram0_READDATAVALID  (ddr_read_readdatavalid),            //                   .readdatavalid
		.f2h_sdram0_READ           (ddr_read_read),                     //                   .read
		.f2h_sdram1_clk            (ddr_write_clock_clk),               //   f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS        (ddr_write_address),                 //    f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT     (ddr_write_burstcount),              //                   .burstcount
		.f2h_sdram1_WAITREQUEST    (ddr_write_waitrequest),             //                   .waitrequest
		.f2h_sdram1_WRITEDATA      (ddr_write_writedata),               //                   .writedata
		.f2h_sdram1_BYTEENABLE     (ddr_write_byteenable),              //                   .byteenable
		.f2h_sdram1_WRITE          (ddr_write_write),                   //                   .write
		.h2f_axi_clk               (user_clock_clk),                    //      h2f_axi_clock.clk
		.h2f_AWID                  (arm_hps_h2f_axi_master_awid),       //     h2f_axi_master.awid
		.h2f_AWADDR                (arm_hps_h2f_axi_master_awaddr),     //                   .awaddr
		.h2f_AWLEN                 (arm_hps_h2f_axi_master_awlen),      //                   .awlen
		.h2f_AWSIZE                (arm_hps_h2f_axi_master_awsize),     //                   .awsize
		.h2f_AWBURST               (arm_hps_h2f_axi_master_awburst),    //                   .awburst
		.h2f_AWLOCK                (arm_hps_h2f_axi_master_awlock),     //                   .awlock
		.h2f_AWCACHE               (arm_hps_h2f_axi_master_awcache),    //                   .awcache
		.h2f_AWPROT                (arm_hps_h2f_axi_master_awprot),     //                   .awprot
		.h2f_AWVALID               (arm_hps_h2f_axi_master_awvalid),    //                   .awvalid
		.h2f_AWREADY               (arm_hps_h2f_axi_master_awready),    //                   .awready
		.h2f_WID                   (arm_hps_h2f_axi_master_wid),        //                   .wid
		.h2f_WDATA                 (arm_hps_h2f_axi_master_wdata),      //                   .wdata
		.h2f_WSTRB                 (arm_hps_h2f_axi_master_wstrb),      //                   .wstrb
		.h2f_WLAST                 (arm_hps_h2f_axi_master_wlast),      //                   .wlast
		.h2f_WVALID                (arm_hps_h2f_axi_master_wvalid),     //                   .wvalid
		.h2f_WREADY                (arm_hps_h2f_axi_master_wready),     //                   .wready
		.h2f_BID                   (arm_hps_h2f_axi_master_bid),        //                   .bid
		.h2f_BRESP                 (arm_hps_h2f_axi_master_bresp),      //                   .bresp
		.h2f_BVALID                (arm_hps_h2f_axi_master_bvalid),     //                   .bvalid
		.h2f_BREADY                (arm_hps_h2f_axi_master_bready),     //                   .bready
		.h2f_ARID                  (arm_hps_h2f_axi_master_arid),       //                   .arid
		.h2f_ARADDR                (arm_hps_h2f_axi_master_araddr),     //                   .araddr
		.h2f_ARLEN                 (arm_hps_h2f_axi_master_arlen),      //                   .arlen
		.h2f_ARSIZE                (arm_hps_h2f_axi_master_arsize),     //                   .arsize
		.h2f_ARBURST               (arm_hps_h2f_axi_master_arburst),    //                   .arburst
		.h2f_ARLOCK                (arm_hps_h2f_axi_master_arlock),     //                   .arlock
		.h2f_ARCACHE               (arm_hps_h2f_axi_master_arcache),    //                   .arcache
		.h2f_ARPROT                (arm_hps_h2f_axi_master_arprot),     //                   .arprot
		.h2f_ARVALID               (arm_hps_h2f_axi_master_arvalid),    //                   .arvalid
		.h2f_ARREADY               (arm_hps_h2f_axi_master_arready),    //                   .arready
		.h2f_RID                   (arm_hps_h2f_axi_master_rid),        //                   .rid
		.h2f_RDATA                 (arm_hps_h2f_axi_master_rdata),      //                   .rdata
		.h2f_RRESP                 (arm_hps_h2f_axi_master_rresp),      //                   .rresp
		.h2f_RLAST                 (arm_hps_h2f_axi_master_rlast),      //                   .rlast
		.h2f_RVALID                (arm_hps_h2f_axi_master_rvalid),     //                   .rvalid
		.h2f_RREADY                (arm_hps_h2f_axi_master_rready),     //                   .rready
		.h2f_lw_axi_clk            (user_clock_clk),                    //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID               (arm_hps_h2f_lw_axi_master_awid),    //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR             (arm_hps_h2f_lw_axi_master_awaddr),  //                   .awaddr
		.h2f_lw_AWLEN              (arm_hps_h2f_lw_axi_master_awlen),   //                   .awlen
		.h2f_lw_AWSIZE             (arm_hps_h2f_lw_axi_master_awsize),  //                   .awsize
		.h2f_lw_AWBURST            (arm_hps_h2f_lw_axi_master_awburst), //                   .awburst
		.h2f_lw_AWLOCK             (arm_hps_h2f_lw_axi_master_awlock),  //                   .awlock
		.h2f_lw_AWCACHE            (arm_hps_h2f_lw_axi_master_awcache), //                   .awcache
		.h2f_lw_AWPROT             (arm_hps_h2f_lw_axi_master_awprot),  //                   .awprot
		.h2f_lw_AWVALID            (arm_hps_h2f_lw_axi_master_awvalid), //                   .awvalid
		.h2f_lw_AWREADY            (arm_hps_h2f_lw_axi_master_awready), //                   .awready
		.h2f_lw_WID                (arm_hps_h2f_lw_axi_master_wid),     //                   .wid
		.h2f_lw_WDATA              (arm_hps_h2f_lw_axi_master_wdata),   //                   .wdata
		.h2f_lw_WSTRB              (arm_hps_h2f_lw_axi_master_wstrb),   //                   .wstrb
		.h2f_lw_WLAST              (arm_hps_h2f_lw_axi_master_wlast),   //                   .wlast
		.h2f_lw_WVALID             (arm_hps_h2f_lw_axi_master_wvalid),  //                   .wvalid
		.h2f_lw_WREADY             (arm_hps_h2f_lw_axi_master_wready),  //                   .wready
		.h2f_lw_BID                (arm_hps_h2f_lw_axi_master_bid),     //                   .bid
		.h2f_lw_BRESP              (arm_hps_h2f_lw_axi_master_bresp),   //                   .bresp
		.h2f_lw_BVALID             (arm_hps_h2f_lw_axi_master_bvalid),  //                   .bvalid
		.h2f_lw_BREADY             (arm_hps_h2f_lw_axi_master_bready),  //                   .bready
		.h2f_lw_ARID               (arm_hps_h2f_lw_axi_master_arid),    //                   .arid
		.h2f_lw_ARADDR             (arm_hps_h2f_lw_axi_master_araddr),  //                   .araddr
		.h2f_lw_ARLEN              (arm_hps_h2f_lw_axi_master_arlen),   //                   .arlen
		.h2f_lw_ARSIZE             (arm_hps_h2f_lw_axi_master_arsize),  //                   .arsize
		.h2f_lw_ARBURST            (arm_hps_h2f_lw_axi_master_arburst), //                   .arburst
		.h2f_lw_ARLOCK             (arm_hps_h2f_lw_axi_master_arlock),  //                   .arlock
		.h2f_lw_ARCACHE            (arm_hps_h2f_lw_axi_master_arcache), //                   .arcache
		.h2f_lw_ARPROT             (arm_hps_h2f_lw_axi_master_arprot),  //                   .arprot
		.h2f_lw_ARVALID            (arm_hps_h2f_lw_axi_master_arvalid), //                   .arvalid
		.h2f_lw_ARREADY            (arm_hps_h2f_lw_axi_master_arready), //                   .arready
		.h2f_lw_RID                (arm_hps_h2f_lw_axi_master_rid),     //                   .rid
		.h2f_lw_RDATA              (arm_hps_h2f_lw_axi_master_rdata),   //                   .rdata
		.h2f_lw_RRESP              (arm_hps_h2f_lw_axi_master_rresp),   //                   .rresp
		.h2f_lw_RLAST              (arm_hps_h2f_lw_axi_master_rlast),   //                   .rlast
		.h2f_lw_RVALID             (arm_hps_h2f_lw_axi_master_rvalid),  //                   .rvalid
		.h2f_lw_RREADY             (arm_hps_h2f_lw_axi_master_rready),  //                   .rready
		.f2h_irq_p0                (arm_hps_f2h_irq0_irq),              //           f2h_irq0.irq
		.f2h_irq_p1                (arm_hps_f2h_irq1_irq)               //           f2h_irq1.irq
	);

	HPSWrapper_baremetal baremetal (
		.clk         (user_clock_clk),                             //   clk1.clk
		.address     (mm_interconnect_0_baremetal_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_baremetal_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_baremetal_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_baremetal_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_baremetal_s1_write),       //       .write
		.readdata    (mm_interconnect_0_baremetal_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_baremetal_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_baremetal_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) ddr_read_rst (
		.reset_in0      (hpsinitreset_user_reset_reset), // reset_in0.reset
		.clk            (ddr_read_clock_clk),            //       clk.clk
		.reset_out      (ddr_read_reset_reset),          // reset_out.reset
		.reset_req      (),                              // (terminated)
		.reset_req_in0  (1'b0),                          // (terminated)
		.reset_in1      (1'b0),                          // (terminated)
		.reset_req_in1  (1'b0),                          // (terminated)
		.reset_in2      (1'b0),                          // (terminated)
		.reset_req_in2  (1'b0),                          // (terminated)
		.reset_in3      (1'b0),                          // (terminated)
		.reset_req_in3  (1'b0),                          // (terminated)
		.reset_in4      (1'b0),                          // (terminated)
		.reset_req_in4  (1'b0),                          // (terminated)
		.reset_in5      (1'b0),                          // (terminated)
		.reset_req_in5  (1'b0),                          // (terminated)
		.reset_in6      (1'b0),                          // (terminated)
		.reset_req_in6  (1'b0),                          // (terminated)
		.reset_in7      (1'b0),                          // (terminated)
		.reset_req_in7  (1'b0),                          // (terminated)
		.reset_in8      (1'b0),                          // (terminated)
		.reset_req_in8  (1'b0),                          // (terminated)
		.reset_in9      (1'b0),                          // (terminated)
		.reset_req_in9  (1'b0),                          // (terminated)
		.reset_in10     (1'b0),                          // (terminated)
		.reset_req_in10 (1'b0),                          // (terminated)
		.reset_in11     (1'b0),                          // (terminated)
		.reset_req_in11 (1'b0),                          // (terminated)
		.reset_in12     (1'b0),                          // (terminated)
		.reset_req_in12 (1'b0),                          // (terminated)
		.reset_in13     (1'b0),                          // (terminated)
		.reset_req_in13 (1'b0),                          // (terminated)
		.reset_in14     (1'b0),                          // (terminated)
		.reset_req_in14 (1'b0),                          // (terminated)
		.reset_in15     (1'b0),                          // (terminated)
		.reset_req_in15 (1'b0)                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) ddr_write_rst (
		.reset_in0      (hpsinitreset_user_reset_reset), // reset_in0.reset
		.clk            (ddr_write_clock_clk),           //       clk.clk
		.reset_out      (ddr_write_reset_reset),         // reset_out.reset
		.reset_req      (),                              // (terminated)
		.reset_req_in0  (1'b0),                          // (terminated)
		.reset_in1      (1'b0),                          // (terminated)
		.reset_req_in1  (1'b0),                          // (terminated)
		.reset_in2      (1'b0),                          // (terminated)
		.reset_req_in2  (1'b0),                          // (terminated)
		.reset_in3      (1'b0),                          // (terminated)
		.reset_req_in3  (1'b0),                          // (terminated)
		.reset_in4      (1'b0),                          // (terminated)
		.reset_req_in4  (1'b0),                          // (terminated)
		.reset_in5      (1'b0),                          // (terminated)
		.reset_req_in5  (1'b0),                          // (terminated)
		.reset_in6      (1'b0),                          // (terminated)
		.reset_req_in6  (1'b0),                          // (terminated)
		.reset_in7      (1'b0),                          // (terminated)
		.reset_req_in7  (1'b0),                          // (terminated)
		.reset_in8      (1'b0),                          // (terminated)
		.reset_req_in8  (1'b0),                          // (terminated)
		.reset_in9      (1'b0),                          // (terminated)
		.reset_req_in9  (1'b0),                          // (terminated)
		.reset_in10     (1'b0),                          // (terminated)
		.reset_req_in10 (1'b0),                          // (terminated)
		.reset_in11     (1'b0),                          // (terminated)
		.reset_req_in11 (1'b0),                          // (terminated)
		.reset_in12     (1'b0),                          // (terminated)
		.reset_req_in12 (1'b0),                          // (terminated)
		.reset_in13     (1'b0),                          // (terminated)
		.reset_req_in13 (1'b0),                          // (terminated)
		.reset_in14     (1'b0),                          // (terminated)
		.reset_req_in14 (1'b0),                          // (terminated)
		.reset_in15     (1'b0),                          // (terminated)
		.reset_req_in15 (1'b0)                           // (terminated)
	);

	HPSWrapper_handshake handshake (
		.clk        (user_clock_clk),                            //                 clk.clk
		.reset_n    (~user_reset_reset),                         //               reset.reset_n
		.address    (mm_interconnect_1_handshake_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_handshake_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_handshake_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_handshake_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_handshake_s1_readdata),   //                    .readdata
		.in_port    (handshake_in_port),                         // external_connection.export
		.out_port   (handshake_out_port),                        //                    .export
		.irq        (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	avmm_reset_hw #(
		.ACTIVE_LOW_OUT (0)
	) hpsinitreset (
		.clock      (user_clock_clk),                                  //      clock.clk
		.reset      (rst_controller_reset_out_reset),                  //      reset.reset
		.chipsel    (mm_interconnect_1_hpsinitreset_slave_chipselect), //      slave.chipselect
		.write      (mm_interconnect_1_hpsinitreset_slave_write),      //           .write
		.writedata  (mm_interconnect_1_hpsinitreset_slave_writedata),  //           .writedata
		.user_reset (hpsinitreset_user_reset_reset)                    // user_reset.reset
	);

	avmm_width_adapter_hw #(
		.MASTER_HAVE_WAITREQ         (0),
		.SLAVE_HAVE_WAITREQ          (0),
		.MASTER_HAVE_READ            (1),
		.SLAVE_HAVE_READ             (1),
		.MASTER_HAVE_CHIPSEL         (1),
		.SLAVE_HAVE_CHIPSEL          (1),
		.MASTER_HAVE_CLOCKEN         (0),
		.SLAVE_HAVE_CLOCKEN          (0),
		.SLAVE_HAS_BYTE_EN           (1),
		.SLAVE_READ_INVERTED         (0),
		.BRIDGE_IS_READONLY          (0),
		.BRIDGE_IS_WRITEONLY         (0),
		.USE_MASTER_BURST_PACKING    (0),
		.PIPELINE_MASTER_WRITE       (0),
		.PIPELINE_MASTER_READ        (0),
		.SLAVE_BURST_MAX             (0),
		.SLAVE_BURST_WIDTH           (1),
		.MASTER_BURST_MAX            (0),
		.MASTER_BURST_WIDTH          (1),
		.MASTER_MEM_SYMBOL_WIDTH     (32),
		.MASTER_MEM_ADDRESS_WIDTH    (14),
		.SLAVE_MEM_SYMBOL_WIDTH      (32),
		.PACKING_FACTOR              (1),
		.ADDR_WIDTH_DIFF             (0),
		.SLAVE_MEM_ADDRESS_WIDTH     (14),
		.SLAVE_MEM_SYM_ADDRESS_WIDTH (14)
	) hps_avmm_master (
		.clock            (user_clock_clk),                                     //  clock.clk
		.reset            (user_reset_reset),                                   //  reset.reset
		.slave_chip_sel   (mm_interconnect_1_hps_avmm_master_slave_chipselect), //  slave.chipselect
		.slave_read       (mm_interconnect_1_hps_avmm_master_slave_read),       //       .read
		.slave_readdata   (mm_interconnect_1_hps_avmm_master_slave_readdata),   //       .readdata
		.slave_writedata  (mm_interconnect_1_hps_avmm_master_slave_writedata),  //       .writedata
		.slave_write      (mm_interconnect_1_hps_avmm_master_slave_write),      //       .write
		.slave_byte_en    (mm_interconnect_1_hps_avmm_master_slave_byteenable), //       .byteenable
		.slave_address    (mm_interconnect_1_hps_avmm_master_slave_address),    //       .address
		.master_chip_sel  (hps_avmm_master_chipselect),                         // master.chipselect
		.master_read      (hps_avmm_master_read),                               //       .read
		.master_readdata  (hps_avmm_master_readdata),                           //       .readdata
		.master_writedata (hps_avmm_master_writedata),                          //       .writedata
		.master_write     (hps_avmm_master_write),                              //       .write
		.master_byte_en   (hps_avmm_master_byteenable),                         //       .byteenable
		.master_address   (hps_avmm_master_address)                             //       .address
	);

	qsys_iface_change_hw #(
		.WIDTH (1)
	) hps_reset (
		.clock  (user_clock_clk),                // conduit_clock.clk
		.reset  (power_on_reset_reset_reset),    // conduit_reset.reset
		.sigIn  (reset_width_overflow_overflow), //       conduit.overflow
		.sigOut (hps_reset_reset_reset)          //         reset.reset_n
	);

	LT24Display #(
		.WIDTH      (240),
		.HEIGHT     (320),
		.CLOCK_FREQ (50000000),
		.XBITS      (8),
		.YBITS      (9)
	) lt24_fpga (
		.clock        (user_clock_clk),                //       clock.clk
		.globalReset  (hpsinitreset_user_reset_reset), // globalReset.reset
		.resetApp     (user_reset_reset),              //    resetApp.reset
		.LT24CS_n     (lt24_display_cs_n),             //     display.cs_n
		.LT24RS       (lt24_display_rs),               //            .rs
		.LT24Rd_n     (lt24_display_rd_n),             //            .rd_n
		.LT24Wr_n     (lt24_display_wr_n),             //            .wr_n
		.LT24Data     (lt24_display_data),             //            .data
		.LT24LCDOn    (lt24_display_on),               //            .on
		.LT24Reset_n  (lt24_display_rst_n),            //            .rst_n
		.pixelReady   (lt24_data_ready),               //        data.ready
		.pixelData    (lt24_data_data),                //            .data
		.pixelWrite   (lt24_data_write),               //            .write
		.xAddr        (lt24_data_xAddr),               //            .xAddr
		.yAddr        (lt24_data_yAddr),               //            .yAddr
		.pixelRawMode (lt24_mode_raw),                 //        mode.raw
		.cmdReady     (lt24_cmd_ready),                //     command.ready
		.cmdData      (lt24_cmd_data),                 //            .data
		.cmdWrite     (lt24_cmd_write),                //            .write
		.cmdDone      (lt24_cmd_done)                  //            .done
	);

	power_on_reset_hw power_on_reset (
		.reset (power_on_reset_reset_reset), // reset.reset
		.clock (user_clock_clk)              // clock.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset50mhz (
		.reset_in0      (~arm_hps_h2f_reset_reset),   // reset_in0.reset
		.reset_in1      (~hps_reset_reset_reset),     // reset_in1.reset
		.reset_in2      (power_on_reset_reset_reset), // reset_in2.reset
		.clk            (user_clock_clk),             //       clk.clk
		.reset_out      (reset50mhz_reset_out_reset), // reset_out.reset
		.reset_req      (),                           // (terminated)
		.reset_req_in0  (1'b0),                       // (terminated)
		.reset_req_in1  (1'b0),                       // (terminated)
		.reset_req_in2  (1'b0),                       // (terminated)
		.reset_in3      (1'b0),                       // (terminated)
		.reset_req_in3  (1'b0),                       // (terminated)
		.reset_in4      (1'b0),                       // (terminated)
		.reset_req_in4  (1'b0),                       // (terminated)
		.reset_in5      (1'b0),                       // (terminated)
		.reset_req_in5  (1'b0),                       // (terminated)
		.reset_in6      (1'b0),                       // (terminated)
		.reset_req_in6  (1'b0),                       // (terminated)
		.reset_in7      (1'b0),                       // (terminated)
		.reset_req_in7  (1'b0),                       // (terminated)
		.reset_in8      (1'b0),                       // (terminated)
		.reset_req_in8  (1'b0),                       // (terminated)
		.reset_in9      (1'b0),                       // (terminated)
		.reset_req_in9  (1'b0),                       // (terminated)
		.reset_in10     (1'b0),                       // (terminated)
		.reset_req_in10 (1'b0),                       // (terminated)
		.reset_in11     (1'b0),                       // (terminated)
		.reset_req_in11 (1'b0),                       // (terminated)
		.reset_in12     (1'b0),                       // (terminated)
		.reset_req_in12 (1'b0),                       // (terminated)
		.reset_in13     (1'b0),                       // (terminated)
		.reset_req_in13 (1'b0),                       // (terminated)
		.reset_in14     (1'b0),                       // (terminated)
		.reset_req_in14 (1'b0),                       // (terminated)
		.reset_in15     (1'b0),                       // (terminated)
		.reset_req_in15 (1'b0)                        // (terminated)
	);

	counter_hw #(
		.AUTO_RESET (0),
		.HAS_ENABLE (0),
		.HAS_ZERO   (0),
		.ZERO_EDGE  (0),
		.WIDTH      (10),
		.INCREMENT  (1),
		.ZERO_VALUE (64'b0000000000000000000000000000000000000000000000000000000000000000),
		.MAX_VALUE  (64'b0000000000000000000000000000000000000000000000000000001111111111),
		.INVERT_MSB (0)
	) reset_width (
		.clock      (user_clock_clk),                //    clock.clk
		.reset      (power_on_reset_reset_reset),    //    reset.reset
		.countValue (),                              //  counter.export
		.overflow   (reset_width_overflow_overflow)  // overflow.overflow
	);

	HPSWrapper_sysid sysid (
		.clock    (user_clock_clk),                                 //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	loanio_uart_hw #(
		.INCLUDE_SYNCHRONISER (1)
	) usb_uart (
		.loan_io_in  (arm_hps_h2f_loan_io_in), // loan_io.in
		.loan_io_oe  (usb_uart_loan_io_oe),    //        .oe
		.loan_io_out (usb_uart_loan_io_out),   //        .out
		.uart_rx     (usb_uart_rx),            //    uart.rx
		.uart_tx     (usb_uart_tx),            //        .tx
		.clock       (user_clock_clk)          //   clock.clk
	);

	HPSWrapper_mm_interconnect_0 mm_interconnect_0 (
		.arm_hps_h2f_axi_master_awid                                        (arm_hps_h2f_axi_master_awid),                //                                       arm_hps_h2f_axi_master.awid
		.arm_hps_h2f_axi_master_awaddr                                      (arm_hps_h2f_axi_master_awaddr),              //                                                             .awaddr
		.arm_hps_h2f_axi_master_awlen                                       (arm_hps_h2f_axi_master_awlen),               //                                                             .awlen
		.arm_hps_h2f_axi_master_awsize                                      (arm_hps_h2f_axi_master_awsize),              //                                                             .awsize
		.arm_hps_h2f_axi_master_awburst                                     (arm_hps_h2f_axi_master_awburst),             //                                                             .awburst
		.arm_hps_h2f_axi_master_awlock                                      (arm_hps_h2f_axi_master_awlock),              //                                                             .awlock
		.arm_hps_h2f_axi_master_awcache                                     (arm_hps_h2f_axi_master_awcache),             //                                                             .awcache
		.arm_hps_h2f_axi_master_awprot                                      (arm_hps_h2f_axi_master_awprot),              //                                                             .awprot
		.arm_hps_h2f_axi_master_awvalid                                     (arm_hps_h2f_axi_master_awvalid),             //                                                             .awvalid
		.arm_hps_h2f_axi_master_awready                                     (arm_hps_h2f_axi_master_awready),             //                                                             .awready
		.arm_hps_h2f_axi_master_wid                                         (arm_hps_h2f_axi_master_wid),                 //                                                             .wid
		.arm_hps_h2f_axi_master_wdata                                       (arm_hps_h2f_axi_master_wdata),               //                                                             .wdata
		.arm_hps_h2f_axi_master_wstrb                                       (arm_hps_h2f_axi_master_wstrb),               //                                                             .wstrb
		.arm_hps_h2f_axi_master_wlast                                       (arm_hps_h2f_axi_master_wlast),               //                                                             .wlast
		.arm_hps_h2f_axi_master_wvalid                                      (arm_hps_h2f_axi_master_wvalid),              //                                                             .wvalid
		.arm_hps_h2f_axi_master_wready                                      (arm_hps_h2f_axi_master_wready),              //                                                             .wready
		.arm_hps_h2f_axi_master_bid                                         (arm_hps_h2f_axi_master_bid),                 //                                                             .bid
		.arm_hps_h2f_axi_master_bresp                                       (arm_hps_h2f_axi_master_bresp),               //                                                             .bresp
		.arm_hps_h2f_axi_master_bvalid                                      (arm_hps_h2f_axi_master_bvalid),              //                                                             .bvalid
		.arm_hps_h2f_axi_master_bready                                      (arm_hps_h2f_axi_master_bready),              //                                                             .bready
		.arm_hps_h2f_axi_master_arid                                        (arm_hps_h2f_axi_master_arid),                //                                                             .arid
		.arm_hps_h2f_axi_master_araddr                                      (arm_hps_h2f_axi_master_araddr),              //                                                             .araddr
		.arm_hps_h2f_axi_master_arlen                                       (arm_hps_h2f_axi_master_arlen),               //                                                             .arlen
		.arm_hps_h2f_axi_master_arsize                                      (arm_hps_h2f_axi_master_arsize),              //                                                             .arsize
		.arm_hps_h2f_axi_master_arburst                                     (arm_hps_h2f_axi_master_arburst),             //                                                             .arburst
		.arm_hps_h2f_axi_master_arlock                                      (arm_hps_h2f_axi_master_arlock),              //                                                             .arlock
		.arm_hps_h2f_axi_master_arcache                                     (arm_hps_h2f_axi_master_arcache),             //                                                             .arcache
		.arm_hps_h2f_axi_master_arprot                                      (arm_hps_h2f_axi_master_arprot),              //                                                             .arprot
		.arm_hps_h2f_axi_master_arvalid                                     (arm_hps_h2f_axi_master_arvalid),             //                                                             .arvalid
		.arm_hps_h2f_axi_master_arready                                     (arm_hps_h2f_axi_master_arready),             //                                                             .arready
		.arm_hps_h2f_axi_master_rid                                         (arm_hps_h2f_axi_master_rid),                 //                                                             .rid
		.arm_hps_h2f_axi_master_rdata                                       (arm_hps_h2f_axi_master_rdata),               //                                                             .rdata
		.arm_hps_h2f_axi_master_rresp                                       (arm_hps_h2f_axi_master_rresp),               //                                                             .rresp
		.arm_hps_h2f_axi_master_rlast                                       (arm_hps_h2f_axi_master_rlast),               //                                                             .rlast
		.arm_hps_h2f_axi_master_rvalid                                      (arm_hps_h2f_axi_master_rvalid),              //                                                             .rvalid
		.arm_hps_h2f_axi_master_rready                                      (arm_hps_h2f_axi_master_rready),              //                                                             .rready
		.clk50mhz_out_clk_clk                                               (user_clock_clk),                             //                                             clk50mhz_out_clk.clk
		.arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),         // arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.baremetal_reset1_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),             //                       baremetal_reset1_reset_bridge_in_reset.reset
		.baremetal_s1_address                                               (mm_interconnect_0_baremetal_s1_address),     //                                                 baremetal_s1.address
		.baremetal_s1_write                                                 (mm_interconnect_0_baremetal_s1_write),       //                                                             .write
		.baremetal_s1_readdata                                              (mm_interconnect_0_baremetal_s1_readdata),    //                                                             .readdata
		.baremetal_s1_writedata                                             (mm_interconnect_0_baremetal_s1_writedata),   //                                                             .writedata
		.baremetal_s1_byteenable                                            (mm_interconnect_0_baremetal_s1_byteenable),  //                                                             .byteenable
		.baremetal_s1_chipselect                                            (mm_interconnect_0_baremetal_s1_chipselect),  //                                                             .chipselect
		.baremetal_s1_clken                                                 (mm_interconnect_0_baremetal_s1_clken),       //                                                             .clken
		.baremetal_s1_debugaccess                                           (mm_interconnect_0_baremetal_s1_debugaccess)  //                                                             .debugaccess
	);

	HPSWrapper_mm_interconnect_1 mm_interconnect_1 (
		.arm_hps_h2f_lw_axi_master_awid                                        (arm_hps_h2f_lw_axi_master_awid),                     //                                       arm_hps_h2f_lw_axi_master.awid
		.arm_hps_h2f_lw_axi_master_awaddr                                      (arm_hps_h2f_lw_axi_master_awaddr),                   //                                                                .awaddr
		.arm_hps_h2f_lw_axi_master_awlen                                       (arm_hps_h2f_lw_axi_master_awlen),                    //                                                                .awlen
		.arm_hps_h2f_lw_axi_master_awsize                                      (arm_hps_h2f_lw_axi_master_awsize),                   //                                                                .awsize
		.arm_hps_h2f_lw_axi_master_awburst                                     (arm_hps_h2f_lw_axi_master_awburst),                  //                                                                .awburst
		.arm_hps_h2f_lw_axi_master_awlock                                      (arm_hps_h2f_lw_axi_master_awlock),                   //                                                                .awlock
		.arm_hps_h2f_lw_axi_master_awcache                                     (arm_hps_h2f_lw_axi_master_awcache),                  //                                                                .awcache
		.arm_hps_h2f_lw_axi_master_awprot                                      (arm_hps_h2f_lw_axi_master_awprot),                   //                                                                .awprot
		.arm_hps_h2f_lw_axi_master_awvalid                                     (arm_hps_h2f_lw_axi_master_awvalid),                  //                                                                .awvalid
		.arm_hps_h2f_lw_axi_master_awready                                     (arm_hps_h2f_lw_axi_master_awready),                  //                                                                .awready
		.arm_hps_h2f_lw_axi_master_wid                                         (arm_hps_h2f_lw_axi_master_wid),                      //                                                                .wid
		.arm_hps_h2f_lw_axi_master_wdata                                       (arm_hps_h2f_lw_axi_master_wdata),                    //                                                                .wdata
		.arm_hps_h2f_lw_axi_master_wstrb                                       (arm_hps_h2f_lw_axi_master_wstrb),                    //                                                                .wstrb
		.arm_hps_h2f_lw_axi_master_wlast                                       (arm_hps_h2f_lw_axi_master_wlast),                    //                                                                .wlast
		.arm_hps_h2f_lw_axi_master_wvalid                                      (arm_hps_h2f_lw_axi_master_wvalid),                   //                                                                .wvalid
		.arm_hps_h2f_lw_axi_master_wready                                      (arm_hps_h2f_lw_axi_master_wready),                   //                                                                .wready
		.arm_hps_h2f_lw_axi_master_bid                                         (arm_hps_h2f_lw_axi_master_bid),                      //                                                                .bid
		.arm_hps_h2f_lw_axi_master_bresp                                       (arm_hps_h2f_lw_axi_master_bresp),                    //                                                                .bresp
		.arm_hps_h2f_lw_axi_master_bvalid                                      (arm_hps_h2f_lw_axi_master_bvalid),                   //                                                                .bvalid
		.arm_hps_h2f_lw_axi_master_bready                                      (arm_hps_h2f_lw_axi_master_bready),                   //                                                                .bready
		.arm_hps_h2f_lw_axi_master_arid                                        (arm_hps_h2f_lw_axi_master_arid),                     //                                                                .arid
		.arm_hps_h2f_lw_axi_master_araddr                                      (arm_hps_h2f_lw_axi_master_araddr),                   //                                                                .araddr
		.arm_hps_h2f_lw_axi_master_arlen                                       (arm_hps_h2f_lw_axi_master_arlen),                    //                                                                .arlen
		.arm_hps_h2f_lw_axi_master_arsize                                      (arm_hps_h2f_lw_axi_master_arsize),                   //                                                                .arsize
		.arm_hps_h2f_lw_axi_master_arburst                                     (arm_hps_h2f_lw_axi_master_arburst),                  //                                                                .arburst
		.arm_hps_h2f_lw_axi_master_arlock                                      (arm_hps_h2f_lw_axi_master_arlock),                   //                                                                .arlock
		.arm_hps_h2f_lw_axi_master_arcache                                     (arm_hps_h2f_lw_axi_master_arcache),                  //                                                                .arcache
		.arm_hps_h2f_lw_axi_master_arprot                                      (arm_hps_h2f_lw_axi_master_arprot),                   //                                                                .arprot
		.arm_hps_h2f_lw_axi_master_arvalid                                     (arm_hps_h2f_lw_axi_master_arvalid),                  //                                                                .arvalid
		.arm_hps_h2f_lw_axi_master_arready                                     (arm_hps_h2f_lw_axi_master_arready),                  //                                                                .arready
		.arm_hps_h2f_lw_axi_master_rid                                         (arm_hps_h2f_lw_axi_master_rid),                      //                                                                .rid
		.arm_hps_h2f_lw_axi_master_rdata                                       (arm_hps_h2f_lw_axi_master_rdata),                    //                                                                .rdata
		.arm_hps_h2f_lw_axi_master_rresp                                       (arm_hps_h2f_lw_axi_master_rresp),                    //                                                                .rresp
		.arm_hps_h2f_lw_axi_master_rlast                                       (arm_hps_h2f_lw_axi_master_rlast),                    //                                                                .rlast
		.arm_hps_h2f_lw_axi_master_rvalid                                      (arm_hps_h2f_lw_axi_master_rvalid),                   //                                                                .rvalid
		.arm_hps_h2f_lw_axi_master_rready                                      (arm_hps_h2f_lw_axi_master_rready),                   //                                                                .rready
		.clk50mhz_out_clk_clk                                                  (user_clock_clk),                                     //                                                clk50mhz_out_clk.clk
		.arm_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                 // arm_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.handshake_reset_reset_bridge_in_reset_reset                           (user_reset_reset),                                   //                           handshake_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                     //                               sysid_reset_reset_bridge_in_reset.reset
		.handshake_s1_address                                                  (mm_interconnect_1_handshake_s1_address),             //                                                    handshake_s1.address
		.handshake_s1_write                                                    (mm_interconnect_1_handshake_s1_write),               //                                                                .write
		.handshake_s1_readdata                                                 (mm_interconnect_1_handshake_s1_readdata),            //                                                                .readdata
		.handshake_s1_writedata                                                (mm_interconnect_1_handshake_s1_writedata),           //                                                                .writedata
		.handshake_s1_chipselect                                               (mm_interconnect_1_handshake_s1_chipselect),          //                                                                .chipselect
		.hps_avmm_master_slave_address                                         (mm_interconnect_1_hps_avmm_master_slave_address),    //                                           hps_avmm_master_slave.address
		.hps_avmm_master_slave_write                                           (mm_interconnect_1_hps_avmm_master_slave_write),      //                                                                .write
		.hps_avmm_master_slave_read                                            (mm_interconnect_1_hps_avmm_master_slave_read),       //                                                                .read
		.hps_avmm_master_slave_readdata                                        (mm_interconnect_1_hps_avmm_master_slave_readdata),   //                                                                .readdata
		.hps_avmm_master_slave_writedata                                       (mm_interconnect_1_hps_avmm_master_slave_writedata),  //                                                                .writedata
		.hps_avmm_master_slave_byteenable                                      (mm_interconnect_1_hps_avmm_master_slave_byteenable), //                                                                .byteenable
		.hps_avmm_master_slave_chipselect                                      (mm_interconnect_1_hps_avmm_master_slave_chipselect), //                                                                .chipselect
		.hpsInitReset_slave_write                                              (mm_interconnect_1_hpsinitreset_slave_write),         //                                              hpsInitReset_slave.write
		.hpsInitReset_slave_writedata                                          (mm_interconnect_1_hpsinitreset_slave_writedata),     //                                                                .writedata
		.hpsInitReset_slave_chipselect                                         (mm_interconnect_1_hpsinitreset_slave_chipselect),    //                                                                .chipselect
		.sysid_control_slave_address                                           (mm_interconnect_1_sysid_control_slave_address),      //                                             sysid_control_slave.address
		.sysid_control_slave_readdata                                          (mm_interconnect_1_sysid_control_slave_readdata)      //                                                                .readdata
	);

	HPSWrapper_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_hps_f2h_irq0_irq)      //    sender.irq
	);

	HPSWrapper_irq_mapper_001 irq_mapper_001 (
		.clk        (),                     //       clk.clk
		.reset      (),                     // clk_reset.reset
		.sender_irq (arm_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset50mhz_reset_out_reset),         // reset_in0.reset
		.clk            (user_clock_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (user_clock_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
